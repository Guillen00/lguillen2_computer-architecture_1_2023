module adder (input [31:0] A,
					input [31:0] B,
					output [31:0] C
	);
	
	//Realiza una suma
	assign C = A + B;
	
endmodule